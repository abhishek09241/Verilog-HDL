`define TRUE  1'b1
`define FALSE 1'b0


// Delays
`define Y2RDELAY 3 // Yellow to Red delay
`define R2YDELAY 2 // Red to Yellow delay


module traffic_signal_control (
    
);
    
endmodule